* C:\Users\DELL\Desktop\LTSPICENETLIST\GPIO_BIDIBUFF_TANVI.asc
M1 from_pad from_pad vdd N009 PMOS
M2 vdd from_pad N012 N010 PMOS
M3 vdd N012 to_core N011 PMOS
M5 N012 from_pad 0 N014 NMOS
M6 to_core N012 0 N015 NMOS
M4 0 from_pad from_pad N013 NMOS
V1 from_pad 0 PULSE(0 2 0 1m 1m 7m 10m)
M7 Vdd Vdd N006 N004 NMOS
M8 Vdd from_int_ckt out_to_pad N005 NMOS
M9 N006 from_int_ckt 0 N007 NMOS
M10 out_to_pad N006 0 N008 NMOS
V2 from_int_ckt 0 PULSE(0 2 0 1m 1m 7m 10m)
M11 N001 N003 0 0 NMOS
M12 Vdd N003 N001 N002 PMOS
V�ENABLE N003 0 PULSE(0 2 0 1m 1m 7m 10m)
.model NMOS NMOS
.model PMOS PMOS
.lib C:\Users\DELL\Documents\LTspiceXVII\lib\cmp\standard.mos
Vdd Vdd 0 DC 3.8
.tran 100m
.backanno
.end
